class monitor
