this is test trail
